class	component;

	virtual	task	build();
	endtask
	virtual	task	reset();
	endtask
	virtual	task	run(int i);
	endtask
	virtual	task	check(int i);
	endtask
	virtual	task	report();
	endtask

endclass

